`timescale 1ns/1ps

module InstructionMemory (Address,Instruction);
input [31:0] Address;
output reg[31:0] Instruction;

always@(*)
    case(Address[10:2])

 9'd0:  Instruction<=32'h08100003;
 9'd1:  Instruction<=32'h08100053;
 9'd2:  Instruction<=32'h081000b7;
 9'd3:  Instruction<=32'h20150001;
 9'd4:  Instruction<=32'h0015af80;
 9'd5:  Instruction<=32'haea00008;
 9'd6:  Instruction<=32'h00004020;
 9'd7:  Instruction<=32'h3c08ffff;
 9'd8:  Instruction<=32'h3c010000;
 9'd9:  Instruction<=32'h3421f52f;
 9'd10:  Instruction<=32'h01014020;
 9'd11:  Instruction<=32'haea80000;
 9'd12:  Instruction<=32'h00004020;
 9'd13:  Instruction<=32'h3c08ffff;
 9'd14:  Instruction<=32'h3c010000;
 9'd15:  Instruction<=32'h3421ffff;
 9'd16:  Instruction<=32'h01014020;
 9'd17:  Instruction<=32'haea80004;
 9'd18:  Instruction<=32'h0c1000b8;
 9'd19:  Instruction<=32'h8c110000;
 9'd20:  Instruction<=32'h2231ffff;
 9'd21:  Instruction<=32'h20100000;
 9'd22:  Instruction<=32'h22100004;
 9'd23:  Instruction<=32'h8eb60014;
 9'd24:  Instruction<=32'h0c10002a;
 9'd25:  Instruction<=32'h8eb70014;
 9'd26:  Instruction<=32'h02f6b822;
 9'd27:  Instruction<=32'h20080003;
 9'd28:  Instruction<=32'haea80008;
 9'd29:  Instruction<=32'h0000a020;
 9'd30:  Instruction<=32'h200e07d0;
 9'd31:  Instruction<=32'h11d40001;
 9'd32:  Instruction<=32'h0810001f;
 9'd33:  Instruction<=32'h0000a020;
 9'd34:  Instruction<=32'h200e07d0;
 9'd35:  Instruction<=32'h8e170000;
 9'd36:  Instruction<=32'h11d40001;
 9'd37:  Instruction<=32'h08100024;
 9'd38:  Instruction<=32'h22100004;
 9'd39:  Instruction<=32'h2231fffc;
 9'd40:  Instruction<=32'h1220015b;
 9'd41:  Instruction<=32'h08100021;
 9'd42:  Instruction<=32'h23bdffec;
 9'd43:  Instruction<=32'hafbf0010;
 9'd44:  Instruction<=32'hafb8000c;
 9'd45:  Instruction<=32'hafaf0008;
 9'd46:  Instruction<=32'hafae0004;
 9'd47:  Instruction<=32'hafad0000;
 9'd48:  Instruction<=32'h00107821;
 9'd49:  Instruction<=32'h0011c021;
 9'd50:  Instruction<=32'h00006821;
 9'd51:  Instruction<=32'h01b8402a;
 9'd52:  Instruction<=32'h11000010;
 9'd53:  Instruction<=32'h21aeffff;
 9'd54:  Instruction<=32'h29c80000;
 9'd55:  Instruction<=32'h1500000b;
 9'd56:  Instruction<=32'h000e4880;
 9'd57:  Instruction<=32'h01e95020;
 9'd58:  Instruction<=32'h8d4b0000;
 9'd59:  Instruction<=32'h8d4c0004;
 9'd60:  Instruction<=32'h018b402a;
 9'd61:  Instruction<=32'h11000005;
 9'd62:  Instruction<=32'h000f8021;
 9'd63:  Instruction<=32'h000e8821;
 9'd64:  Instruction<=32'h0c10004c;
 9'd65:  Instruction<=32'h21ceffff;
 9'd66:  Instruction<=32'h08100036;
 9'd67:  Instruction<=32'h21ad0001;
 9'd68:  Instruction<=32'h08100033;
 9'd69:  Instruction<=32'h8fad0000;
 9'd70:  Instruction<=32'h8fae0004;
 9'd71:  Instruction<=32'h8faf0008;
 9'd72:  Instruction<=32'h8fb8000c;
 9'd73:  Instruction<=32'h8fbf0010;
 9'd74:  Instruction<=32'h23bd0014;
 9'd75:  Instruction<=32'h03e00008;
 9'd76:  Instruction<=32'h00114880;
 9'd77:  Instruction<=32'h02094820;
 9'd78:  Instruction<=32'h8d280000;
 9'd79:  Instruction<=32'h8d2a0004;
 9'd80:  Instruction<=32'had2a0000;
 9'd81:  Instruction<=32'had280004;
 9'd82:  Instruction<=32'h03e00008;
 9'd83:  Instruction<=32'haea00008;
 9'd84:  Instruction<=32'h22940001;
 9'd85:  Instruction<=32'h20120003;
 9'd86:  Instruction<=32'h02929824;
 9'd87:  Instruction<=32'h200a000f;
 9'd88:  Instruction<=32'h20080000;
 9'd89:  Instruction<=32'h12680006;
 9'd90:  Instruction<=32'h20080001;
 9'd91:  Instruction<=32'h12680007;
 9'd92:  Instruction<=32'h20080002;
 9'd93:  Instruction<=32'h1268000a;
 9'd94:  Instruction<=32'h20080003;
 9'd95:  Instruction<=32'h1268000d;
 9'd96:  Instruction<=32'h02ea4824;
 9'd97:  Instruction<=32'h200c000e;
 9'd98:  Instruction<=32'h08100072;
 9'd99:  Instruction<=32'h000a5100;
 9'd100:  Instruction<=32'h02ea4824;
 9'd101:  Instruction<=32'h00094902;
 9'd102:  Instruction<=32'h200c000d;
 9'd103:  Instruction<=32'h08100072;
 9'd104:  Instruction<=32'h000a5200;
 9'd105:  Instruction<=32'h02ea4824;
 9'd106:  Instruction<=32'h00094a02;
 9'd107:  Instruction<=32'h200c000b;
 9'd108:  Instruction<=32'h08100072;
 9'd109:  Instruction<=32'h000a5300;
 9'd110:  Instruction<=32'h02ea4824;
 9'd111:  Instruction<=32'h00094b02;
 9'd112:  Instruction<=32'h200c0007;
 9'd113:  Instruction<=32'h08100072;
 9'd114:  Instruction<=32'h000c6200;
 9'd115:  Instruction<=32'h200b0000;
 9'd116:  Instruction<=32'h112b001e;
 9'd117:  Instruction<=32'h200b0001;
 9'd118:  Instruction<=32'h112b001e;
 9'd119:  Instruction<=32'h200b0002;
 9'd120:  Instruction<=32'h112b001e;
 9'd121:  Instruction<=32'h200b0003;
 9'd122:  Instruction<=32'h112b001e;
 9'd123:  Instruction<=32'h200b0004;
 9'd124:  Instruction<=32'h112b001e;
 9'd125:  Instruction<=32'h200b0005;
 9'd126:  Instruction<=32'h112b001e;
 9'd127:  Instruction<=32'h200b0006;
 9'd128:  Instruction<=32'h112b001e;
 9'd129:  Instruction<=32'h200b0007;
 9'd130:  Instruction<=32'h112b001e;
 9'd131:  Instruction<=32'h200b0008;
 9'd132:  Instruction<=32'h112b001e;
 9'd133:  Instruction<=32'h200b0009;
 9'd134:  Instruction<=32'h112b001e;
 9'd135:  Instruction<=32'h200b000a;
 9'd136:  Instruction<=32'h112b001e;
 9'd137:  Instruction<=32'h200b000b;
 9'd138:  Instruction<=32'h112b001e;
 9'd139:  Instruction<=32'h200b000c;
 9'd140:  Instruction<=32'h112b001e;
 9'd141:  Instruction<=32'h200b000d;
 9'd142:  Instruction<=32'h112b001e;
 9'd143:  Instruction<=32'h200b000e;
 9'd144:  Instruction<=32'h112b001e;
 9'd145:  Instruction<=32'h200b000f;
 9'd146:  Instruction<=32'h112b001e;
 9'd147:  Instruction<=32'h218d0040;
 9'd148:  Instruction<=32'h081000b3;
 9'd149:  Instruction<=32'h218d0079;
 9'd150:  Instruction<=32'h081000b3;
 9'd151:  Instruction<=32'h218d0024;
 9'd152:  Instruction<=32'h081000b3;
 9'd153:  Instruction<=32'h218d0030;
 9'd154:  Instruction<=32'h081000b3;
 9'd155:  Instruction<=32'h218d0019;
 9'd156:  Instruction<=32'h081000b3;
 9'd157:  Instruction<=32'h218d0012;
 9'd158:  Instruction<=32'h081000b3;
 9'd159:  Instruction<=32'h218d0002;
 9'd160:  Instruction<=32'h081000b3;
 9'd161:  Instruction<=32'h218d0078;
 9'd162:  Instruction<=32'h081000b3;
 9'd163:  Instruction<=32'h218d0000;
 9'd164:  Instruction<=32'h081000b3;
 9'd165:  Instruction<=32'h218d0010;
 9'd166:  Instruction<=32'h081000b3;
 9'd167:  Instruction<=32'h218d0008;
 9'd168:  Instruction<=32'h081000b3;
 9'd169:  Instruction<=32'h218d0003;
 9'd170:  Instruction<=32'h081000b3;
 9'd171:  Instruction<=32'h218d0046;
 9'd172:  Instruction<=32'h081000b3;
 9'd173:  Instruction<=32'h218d0021;
 9'd174:  Instruction<=32'h081000b3;
 9'd175:  Instruction<=32'h218d0006;
 9'd176:  Instruction<=32'h081000b3;
 9'd177:  Instruction<=32'h218d000e;
 9'd178:  Instruction<=32'h081000b3;
 9'd179:  Instruction<=32'haead0010;
 9'd180:  Instruction<=32'h20080003;
 9'd181:  Instruction<=32'haea80008;
 9'd182:  Instruction<=32'h03400008;
 9'd183:  Instruction<=32'h081000b7;
 9'd184:  Instruction<=32'h20090000;
 9'd185:  Instruction<=32'h20080064;
 9'd186:  Instruction<=32'had280000;
 9'd187:  Instruction<=32'h200801d4;
 9'd188:  Instruction<=32'had280004;
 9'd189:  Instruction<=32'h200800e9;
 9'd190:  Instruction<=32'had280008;
 9'd191:  Instruction<=32'h20080151;
 9'd192:  Instruction<=32'had28000c;
 9'd193:  Instruction<=32'h200801f2;
 9'd194:  Instruction<=32'had280010;
 9'd195:  Instruction<=32'h200800ad;
 9'd196:  Instruction<=32'had280014;
 9'd197:  Instruction<=32'h200802d2;
 9'd198:  Instruction<=32'had280018;
 9'd199:  Instruction<=32'h200801dc;
 9'd200:  Instruction<=32'had28001c;
 9'd201:  Instruction<=32'h20080163;
 9'd202:  Instruction<=32'had280020;
 9'd203:  Instruction<=32'h20080060;
 9'd204:  Instruction<=32'had280024;
 9'd205:  Instruction<=32'h200801c8;
 9'd206:  Instruction<=32'had280028;
 9'd207:  Instruction<=32'h200802bf;
 9'd208:  Instruction<=32'had28002c;
 9'd209:  Instruction<=32'h20080082;
 9'd210:  Instruction<=32'had280030;
 9'd211:  Instruction<=32'h2008011c;
 9'd212:  Instruction<=32'had280034;
 9'd213:  Instruction<=32'h2008033d;
 9'd214:  Instruction<=32'had280038;
 9'd215:  Instruction<=32'h200803c7;
 9'd216:  Instruction<=32'had28003c;
 9'd217:  Instruction<=32'h200801e9;
 9'd218:  Instruction<=32'had280040;
 9'd219:  Instruction<=32'h200803a6;
 9'd220:  Instruction<=32'had280044;
 9'd221:  Instruction<=32'h200803e4;
 9'd222:  Instruction<=32'had280048;
 9'd223:  Instruction<=32'h20080189;
 9'd224:  Instruction<=32'had28004c;
 9'd225:  Instruction<=32'h2008002f;
 9'd226:  Instruction<=32'had280050;
 9'd227:  Instruction<=32'h20080366;
 9'd228:  Instruction<=32'had280054;
 9'd229:  Instruction<=32'h2008025f;
 9'd230:  Instruction<=32'had280058;
 9'd231:  Instruction<=32'h20080393;
 9'd232:  Instruction<=32'had28005c;
 9'd233:  Instruction<=32'h2008008f;
 9'd234:  Instruction<=32'had280060;
 9'd235:  Instruction<=32'h2008012a;
 9'd236:  Instruction<=32'had280064;
 9'd237:  Instruction<=32'h20080181;
 9'd238:  Instruction<=32'had280068;
 9'd239:  Instruction<=32'h200801a5;
 9'd240:  Instruction<=32'had28006c;
 9'd241:  Instruction<=32'h200802d7;
 9'd242:  Instruction<=32'had280070;
 9'd243:  Instruction<=32'h200802c5;
 9'd244:  Instruction<=32'had280074;
 9'd245:  Instruction<=32'h20080059;
 9'd246:  Instruction<=32'had280078;
 9'd247:  Instruction<=32'h200801e4;
 9'd248:  Instruction<=32'had28007c;
 9'd249:  Instruction<=32'h200802cd;
 9'd250:  Instruction<=32'had280080;
 9'd251:  Instruction<=32'h20080304;
 9'd252:  Instruction<=32'had280084;
 9'd253:  Instruction<=32'h20080251;
 9'd254:  Instruction<=32'had280088;
 9'd255:  Instruction<=32'h20080331;
 9'd256:  Instruction<=32'had28008c;
 9'd257:  Instruction<=32'h20080391;
 9'd258:  Instruction<=32'had280090;
 9'd259:  Instruction<=32'h2008029d;
 9'd260:  Instruction<=32'had280094;
 9'd261:  Instruction<=32'h2008012c;
 9'd262:  Instruction<=32'had280098;
 9'd263:  Instruction<=32'h20080025;
 9'd264:  Instruction<=32'had28009c;
 9'd265:  Instruction<=32'h2008037f;
 9'd266:  Instruction<=32'had2800a0;
 9'd267:  Instruction<=32'h2008025c;
 9'd268:  Instruction<=32'had2800a4;
 9'd269:  Instruction<=32'h20080200;
 9'd270:  Instruction<=32'had2800a8;
 9'd271:  Instruction<=32'h2008007b;
 9'd272:  Instruction<=32'had2800ac;
 9'd273:  Instruction<=32'h2008014d;
 9'd274:  Instruction<=32'had2800b0;
 9'd275:  Instruction<=32'h2008028a;
 9'd276:  Instruction<=32'had2800b4;
 9'd277:  Instruction<=32'h20080270;
 9'd278:  Instruction<=32'had2800b8;
 9'd279:  Instruction<=32'h2008008b;
 9'd280:  Instruction<=32'had2800bc;
 9'd281:  Instruction<=32'h200802e9;
 9'd282:  Instruction<=32'had2800c0;
 9'd283:  Instruction<=32'h200800fb;
 9'd284:  Instruction<=32'had2800c4;
 9'd285:  Instruction<=32'h200800f6;
 9'd286:  Instruction<=32'had2800c8;
 9'd287:  Instruction<=32'h2008021a;
 9'd288:  Instruction<=32'had2800cc;
 9'd289:  Instruction<=32'h20080285;
 9'd290:  Instruction<=32'had2800d0;
 9'd291:  Instruction<=32'h20080297;
 9'd292:  Instruction<=32'had2800d4;
 9'd293:  Instruction<=32'h200802f6;
 9'd294:  Instruction<=32'had2800d8;
 9'd295:  Instruction<=32'h2008008a;
 9'd296:  Instruction<=32'had2800dc;
 9'd297:  Instruction<=32'h2008035d;
 9'd298:  Instruction<=32'had2800e0;
 9'd299:  Instruction<=32'h2008007c;
 9'd300:  Instruction<=32'had2800e4;
 9'd301:  Instruction<=32'h200803ae;
 9'd302:  Instruction<=32'had2800e8;
 9'd303:  Instruction<=32'h200800e6;
 9'd304:  Instruction<=32'had2800ec;
 9'd305:  Instruction<=32'h20080024;
 9'd306:  Instruction<=32'had2800f0;
 9'd307:  Instruction<=32'h2008013d;
 9'd308:  Instruction<=32'had2800f4;
 9'd309:  Instruction<=32'h200803d2;
 9'd310:  Instruction<=32'had2800f8;
 9'd311:  Instruction<=32'h200800bf;
 9'd312:  Instruction<=32'had2800fc;
 9'd313:  Instruction<=32'h2008006b;
 9'd314:  Instruction<=32'had280100;
 9'd315:  Instruction<=32'h20080121;
 9'd316:  Instruction<=32'had280104;
 9'd317:  Instruction<=32'h20080283;
 9'd318:  Instruction<=32'had280108;
 9'd319:  Instruction<=32'h200803af;
 9'd320:  Instruction<=32'had28010c;
 9'd321:  Instruction<=32'h2008002a;
 9'd322:  Instruction<=32'had280110;
 9'd323:  Instruction<=32'h200801bf;
 9'd324:  Instruction<=32'had280114;
 9'd325:  Instruction<=32'h20080372;
 9'd326:  Instruction<=32'had280118;
 9'd327:  Instruction<=32'h20080109;
 9'd328:  Instruction<=32'had28011c;
 9'd329:  Instruction<=32'h20080326;
 9'd330:  Instruction<=32'had280120;
 9'd331:  Instruction<=32'h2008037b;
 9'd332:  Instruction<=32'had280124;
 9'd333:  Instruction<=32'h20080173;
 9'd334:  Instruction<=32'had280128;
 9'd335:  Instruction<=32'h2008015f;
 9'd336:  Instruction<=32'had28012c;
 9'd337:  Instruction<=32'h2008021c;
 9'd338:  Instruction<=32'had280130;
 9'd339:  Instruction<=32'h20080066;
 9'd340:  Instruction<=32'had280134;
 9'd341:  Instruction<=32'h20080047;
 9'd342:  Instruction<=32'had280138;
 9'd343:  Instruction<=32'h2008018a;
 9'd344:  Instruction<=32'had28013c;
 9'd345:  Instruction<=32'h20080225;
 9'd346:  Instruction<=32'had280140;
 9'd347:  Instruction<=32'h2008027f;
 9'd348:  Instruction<=32'had280144;
 9'd349:  Instruction<=32'h20080269;
 9'd350:  Instruction<=32'had280148;
 9'd351:  Instruction<=32'h20080007;
 9'd352:  Instruction<=32'had28014c;
 9'd353:  Instruction<=32'h200803bb;
 9'd354:  Instruction<=32'had280150;
 9'd355:  Instruction<=32'h200802f5;
 9'd356:  Instruction<=32'had280154;
 9'd357:  Instruction<=32'h20080349;
 9'd358:  Instruction<=32'had280158;
 9'd359:  Instruction<=32'h200803a4;
 9'd360:  Instruction<=32'had28015c;
 9'd361:  Instruction<=32'h20080167;
 9'd362:  Instruction<=32'had280160;
 9'd363:  Instruction<=32'h200803c7;
 9'd364:  Instruction<=32'had280164;
 9'd365:  Instruction<=32'h200801b8;
 9'd366:  Instruction<=32'had280168;
 9'd367:  Instruction<=32'h200803b1;
 9'd368:  Instruction<=32'had28016c;
 9'd369:  Instruction<=32'h200800d1;
 9'd370:  Instruction<=32'had280170;
 9'd371:  Instruction<=32'h20080270;
 9'd372:  Instruction<=32'had280174;
 9'd373:  Instruction<=32'h20080181;
 9'd374:  Instruction<=32'had280178;
 9'd375:  Instruction<=32'h2008021b;
 9'd376:  Instruction<=32'had28017c;
 9'd377:  Instruction<=32'h2008021a;
 9'd378:  Instruction<=32'had280180;
 9'd379:  Instruction<=32'h2008038f;
 9'd380:  Instruction<=32'had280184;
 9'd381:  Instruction<=32'h2008003a;
 9'd382:  Instruction<=32'had280188;
 9'd383:  Instruction<=32'h200803a2;
 9'd384:  Instruction<=32'had28018c;
 9'd385:  Instruction<=32'h2008023c;
 9'd386:  Instruction<=32'had280190;
 9'd387:  Instruction<=32'h03e00008;
 
 default: Instruction<=32'b00000000;

    endcase  
endmodule